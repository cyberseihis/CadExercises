
module div (dig1, dig2, res);
  input [3:0] dig1, dig2;
  output [3:0] res;
  assign res = (dig1 == 4'd0 && dig2 == 4'd0) ? 4'd0 :
(dig1 == 4'd0 && dig2 == 4'd1) ? 4'd0 :
(dig1 == 4'd0 && dig2 == 4'd2) ? 4'd0 :
(dig1 == 4'd0 && dig2 == 4'd3) ? 4'd0 :
(dig1 == 4'd0 && dig2 == 4'd4) ? 4'd0 :
(dig1 == 4'd0 && dig2 == 4'd5) ? 4'd0 :
(dig1 == 4'd0 && dig2 == 4'd6) ? 4'd0 :
(dig1 == 4'd0 && dig2 == 4'd7) ? 4'd0 :
(dig1 == 4'd0 && dig2 == 4'd8) ? 4'd0 :
(dig1 == 4'd0 && dig2 == 4'd9) ? 4'd0 :
(dig1 == 4'd1 && dig2 == 4'd0) ? 4'd0 :
(dig1 == 4'd1 && dig2 == 4'd1) ? 4'd1 :
(dig1 == 4'd1 && dig2 == 4'd2) ? 4'd0 :
(dig1 == 4'd1 && dig2 == 4'd3) ? 4'd0 :
(dig1 == 4'd1 && dig2 == 4'd4) ? 4'd0 :
(dig1 == 4'd1 && dig2 == 4'd5) ? 4'd0 :
(dig1 == 4'd1 && dig2 == 4'd6) ? 4'd0 :
(dig1 == 4'd1 && dig2 == 4'd7) ? 4'd0 :
(dig1 == 4'd1 && dig2 == 4'd8) ? 4'd0 :
(dig1 == 4'd1 && dig2 == 4'd9) ? 4'd0 :
(dig1 == 4'd2 && dig2 == 4'd0) ? 4'd0 :
(dig1 == 4'd2 && dig2 == 4'd1) ? 4'd2 :
(dig1 == 4'd2 && dig2 == 4'd2) ? 4'd1 :
(dig1 == 4'd2 && dig2 == 4'd3) ? 4'd0 :
(dig1 == 4'd2 && dig2 == 4'd4) ? 4'd0 :
(dig1 == 4'd2 && dig2 == 4'd5) ? 4'd0 :
(dig1 == 4'd2 && dig2 == 4'd6) ? 4'd0 :
(dig1 == 4'd2 && dig2 == 4'd7) ? 4'd0 :
(dig1 == 4'd2 && dig2 == 4'd8) ? 4'd0 :
(dig1 == 4'd2 && dig2 == 4'd9) ? 4'd0 :
(dig1 == 4'd3 && dig2 == 4'd0) ? 4'd0 :
(dig1 == 4'd3 && dig2 == 4'd1) ? 4'd3 :
(dig1 == 4'd3 && dig2 == 4'd2) ? 4'd1 :
(dig1 == 4'd3 && dig2 == 4'd3) ? 4'd1 :
(dig1 == 4'd3 && dig2 == 4'd4) ? 4'd0 :
(dig1 == 4'd3 && dig2 == 4'd5) ? 4'd0 :
(dig1 == 4'd3 && dig2 == 4'd6) ? 4'd0 :
(dig1 == 4'd3 && dig2 == 4'd7) ? 4'd0 :
(dig1 == 4'd3 && dig2 == 4'd8) ? 4'd0 :
(dig1 == 4'd3 && dig2 == 4'd9) ? 4'd0 :
(dig1 == 4'd4 && dig2 == 4'd0) ? 4'd0 :
(dig1 == 4'd4 && dig2 == 4'd1) ? 4'd4 :
(dig1 == 4'd4 && dig2 == 4'd2) ? 4'd2 :
(dig1 == 4'd4 && dig2 == 4'd3) ? 4'd1 :
(dig1 == 4'd4 && dig2 == 4'd4) ? 4'd1 :
(dig1 == 4'd4 && dig2 == 4'd5) ? 4'd0 :
(dig1 == 4'd4 && dig2 == 4'd6) ? 4'd0 :
(dig1 == 4'd4 && dig2 == 4'd7) ? 4'd0 :
(dig1 == 4'd4 && dig2 == 4'd8) ? 4'd0 :
(dig1 == 4'd4 && dig2 == 4'd9) ? 4'd0 :
(dig1 == 4'd5 && dig2 == 4'd0) ? 4'd0 :
(dig1 == 4'd5 && dig2 == 4'd1) ? 4'd5 :
(dig1 == 4'd5 && dig2 == 4'd2) ? 4'd2 :
(dig1 == 4'd5 && dig2 == 4'd3) ? 4'd1 :
(dig1 == 4'd5 && dig2 == 4'd4) ? 4'd1 :
(dig1 == 4'd5 && dig2 == 4'd5) ? 4'd1 :
(dig1 == 4'd5 && dig2 == 4'd6) ? 4'd0 :
(dig1 == 4'd5 && dig2 == 4'd7) ? 4'd0 :
(dig1 == 4'd5 && dig2 == 4'd8) ? 4'd0 :
(dig1 == 4'd5 && dig2 == 4'd9) ? 4'd0 :
(dig1 == 4'd6 && dig2 == 4'd0) ? 4'd0 :
(dig1 == 4'd6 && dig2 == 4'd1) ? 4'd6 :
(dig1 == 4'd6 && dig2 == 4'd2) ? 4'd3 :
(dig1 == 4'd6 && dig2 == 4'd3) ? 4'd2 :
(dig1 == 4'd6 && dig2 == 4'd4) ? 4'd1 :
(dig1 == 4'd6 && dig2 == 4'd5) ? 4'd1 :
(dig1 == 4'd6 && dig2 == 4'd6) ? 4'd1 :
(dig1 == 4'd6 && dig2 == 4'd7) ? 4'd0 :
(dig1 == 4'd6 && dig2 == 4'd8) ? 4'd0 :
(dig1 == 4'd6 && dig2 == 4'd9) ? 4'd0 :
(dig1 == 4'd7 && dig2 == 4'd0) ? 4'd0 :
(dig1 == 4'd7 && dig2 == 4'd1) ? 4'd7 :
(dig1 == 4'd7 && dig2 == 4'd2) ? 4'd3 :
(dig1 == 4'd7 && dig2 == 4'd3) ? 4'd2 :
(dig1 == 4'd7 && dig2 == 4'd4) ? 4'd1 :
(dig1 == 4'd7 && dig2 == 4'd5) ? 4'd1 :
(dig1 == 4'd7 && dig2 == 4'd6) ? 4'd1 :
(dig1 == 4'd7 && dig2 == 4'd7) ? 4'd1 :
(dig1 == 4'd7 && dig2 == 4'd8) ? 4'd0 :
(dig1 == 4'd7 && dig2 == 4'd9) ? 4'd0 :
(dig1 == 4'd8 && dig2 == 4'd0) ? 4'd0 :
(dig1 == 4'd8 && dig2 == 4'd1) ? 4'd8 :
(dig1 == 4'd8 && dig2 == 4'd2) ? 4'd4 :
(dig1 == 4'd8 && dig2 == 4'd3) ? 4'd2 :
(dig1 == 4'd8 && dig2 == 4'd4) ? 4'd2 :
(dig1 == 4'd8 && dig2 == 4'd5) ? 4'd1 :
(dig1 == 4'd8 && dig2 == 4'd6) ? 4'd1 :
(dig1 == 4'd8 && dig2 == 4'd7) ? 4'd1 :
(dig1 == 4'd8 && dig2 == 4'd8) ? 4'd1 :
(dig1 == 4'd8 && dig2 == 4'd9) ? 4'd0 :
(dig1 == 4'd9 && dig2 == 4'd0) ? 4'd0 :
(dig1 == 4'd9 && dig2 == 4'd1) ? 4'd9 :
(dig1 == 4'd9 && dig2 == 4'd2) ? 4'd4 :
(dig1 == 4'd9 && dig2 == 4'd3) ? 4'd3 :
(dig1 == 4'd9 && dig2 == 4'd4) ? 4'd2 :
(dig1 == 4'd9 && dig2 == 4'd5) ? 4'd1 :
(dig1 == 4'd9 && dig2 == 4'd6) ? 4'd1 :
(dig1 == 4'd9 && dig2 == 4'd7) ? 4'd1 :
(dig1 == 4'd9 && dig2 == 4'd8) ? 4'd1 :
(dig1 == 4'd9 && dig2 == 4'd9) ? 4'd1 :0;
endmodule